i am in first
