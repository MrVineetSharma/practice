hello i am in second file
